library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity morseDecoder is
	port ( morse: in std_logic_vector (7 downto 0);
			sevenSegment: out std_logic_vector (6 downto 0);
		);
end morseDecoder;
 
architecture arch of morseDecoder is
 
begin
	sevenSegment(0) <= 
	(morse(7) and not morse(6) and not morse(2) and morse(1) and not morse(0))
	or (not morse(7) and not morse(2) and not morse(1) and morse(0))
	or (not morse(7) and morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0))
	or (not morse(7) and morse(6) and morse(5) and not morse(2) and morse(1) and morse(0))
	or (not morse(7) and not morse(6) and not morse(2) and morse(1) and not morse(0))
	or (morse(7) and morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0))
	or (morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0))
	or (morse(7) and morse(6) and not morse(2) and morse(1) and not morse(0))
	or (not morse(7) and morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0))
	or (morse(7) and not morse(6) and morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0))
	or (not morse(7) and not morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0))
	or (morse(7) and morse(6) and morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0))
	or (morse(7) and morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0))
	or (not morse(7) and not morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0))
	or (not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(3) and morse(2) and not morse(1) and morse(0))
	or (not morse(7) and not morse(6) and not morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0))
	or (not morse(7) and not morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0))
	or (not morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0))
	or (morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0));

	sevenSegment(1) <= (and morse(7) and not morse(6) and not morse(2) and morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and not morse(6) and morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0));
	sevenSegment(2) <= (and morse(7) and not morse(6) and not morse(2) and morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(2) and morse(1) and not morse(0)) or (and not morse(7) and morse(6) and not morse(2) and morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and not morse(6) and morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0));
	sevenSegment(3) <= (and morse(7) and not morse(6) and not morse(2) and morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and not morse(2) and not morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and not morse(2) and not morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0));
	sevenSegment(4) <= (and morse(7) and not morse(6) and not morse(2) and morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and not morse(2) and not morse(1) and morse(0)) or (and not morse(7) and morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and not morse(2) and morse(1) and not morse(0)) or (and morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and not morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and not morse(2) and morse(1) and not morse(0)) or (and not morse(7) and morse(6) and not morse(2) and morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and not morse(2) and not morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0));
	sevenSegment(5) <= (and not morse(7) and not morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(2) and not morse(1) and morse(0)) or (and not morse(7) and morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and not morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and not morse(6) and morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and not morse(2) and not morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0))
	sevenSegment(6) <= (and morse(7) and not morse(6) and not morse(2) and morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and not morse(2) and not morse(1) and morse(0)) or (and not morse(7) and morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and not morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(2) and morse(1) and not morse(0)) or (and not morse(7) and morse(6) and not morse(2) and morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(2) and morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and not morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and not morse(6) and morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and not morse(7) and morse(6) and not morse(5) and not morse(2) and morse(1) and morse(0)) or (and morse(7) and not morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(5) and morse(4) and morse(2) and not morse(1) and not morse(0)) or (and morse(7) and morse(6) and morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and morse(7) and not morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and not morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and not morse(5) and not morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and not morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0)) or (and not morse(7) and morse(6) and morse(5) and morse(4) and morse(3) and morse(2) and not morse(1) and morse(0))
end arch;